##
##  Automaticly created by Ofir Even-chen and Yogev Laks Script
####
##  Automaticly created by Ofir Even-chen and Yogev Laks Script
##

VERSION 5.6 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MACRO CDK_R256X16
  CLASS BLOCK ;
  SIZE X_VALUE_SWITCH_LATER BY Y_VALUE_SWITCH_LATER ;
  FOREIGN CDK_R256X16 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN ADDRESS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 12.0 47.0 12.66 47.66 ;
      LAYER Metal6 ;
	RECT 12.0 47.0 12.66 47.66 ;
      LAYER Metal3 ;
	RECT 12.0 47.0 12.66 47.66 ;
      LAYER Metal4 ;
	RECT 12.0 47.0 12.66 47.66 ;
    END
  END ADDRESS[5]
  PIN ADDRESS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 12.0 40.0 12.66 40.66 ;
      LAYER Metal6 ;
	RECT 12.0 40.0 12.66 40.66 ;
      LAYER Metal3 ;
	RECT 12.0 40.0 12.66 40.66 ;
      LAYER Metal4 ;
	RECT 12.0 40.0 12.66 40.66 ;
    END
  END ADDRESS[4]
  PIN ADDRESS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 12.0 33.0 12.66 33.66 ;
      LAYER Metal6 ;
	RECT 12.0 33.0 12.66 33.66 ;
      LAYER Metal3 ;
	RECT 12.0 33.0 12.66 33.66 ;
      LAYER Metal4 ;
	RECT 12.0 33.0 12.66 33.66 ;
    END
  END ADDRESS[3]
  PIN ADDRESS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 12.0 26.0 12.66 26.66 ;
      LAYER Metal6 ;
	RECT 12.0 26.0 12.66 26.66 ;
      LAYER Metal3 ;
	RECT 12.0 26.0 12.66 26.66 ;
      LAYER Metal4 ;
	RECT 12.0 26.0 12.66 26.66 ;
    END
  END ADDRESS[2]
  PIN ADDRESS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 12.0 19.0 12.66 19.66 ;
      LAYER Metal6 ;
	RECT 12.0 19.0 12.66 19.66 ;
      LAYER Metal3 ;
	RECT 12.0 19.0 12.66 19.66 ;
      LAYER Metal4 ;
	RECT 12.0 19.0 12.66 19.66 ;
    END
  END ADDRESS[1]
  PIN ADDRESS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 12.0 12.0 12.66 12.66 ;
      LAYER Metal6 ;
	RECT 12.0 12.0 12.66 12.66 ;
      LAYER Metal3 ;
	RECT 12.0 12.0 12.66 12.66 ;
      LAYER Metal4 ;
	RECT 12.0 12.0 12.66 12.66 ;
    END
  END ADDRESS[0]
  PIN DATA_IN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 26.66 19.66 27.32 20.32 ;
      LAYER Metal6 ;
	RECT 26.66 19.66 27.32 20.32 ;
      LAYER Metal3 ;
	RECT 26.66 19.66 27.32 20.32 ;
      LAYER Metal4 ;
	RECT 26.66 19.66 27.32 20.32 ;
    END
  END DATA_IN[1]
  PIN DATA_IN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 19.66 19.66 20.32 20.32 ;
      LAYER Metal6 ;
	RECT 19.66 19.66 20.32 20.32 ;
      LAYER Metal3 ;
	RECT 19.66 19.66 20.32 20.32 ;
      LAYER Metal4 ;
	RECT 19.66 19.66 20.32 20.32 ;
    END
  END DATA_IN[0]
  PIN DATA_OUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 34.32 27.32 34.98 27.98 ;
      LAYER Metal6 ;
	RECT 34.32 27.32 34.98 27.98 ;
      LAYER Metal3 ;
	RECT 34.32 27.32 34.98 27.98 ;
      LAYER Metal4 ;
	RECT 34.32 27.32 34.98 27.98 ;
    END
  END DATA_OUT[1]
  PIN DATA_OUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 27.32 27.32 27.98 27.98 ;
      LAYER Metal6 ;
	RECT 27.32 27.32 27.98 27.98 ;
      LAYER Metal3 ;
	RECT 27.32 27.32 27.98 27.98 ;
      LAYER Metal4 ;
	RECT 27.32 27.32 27.98 27.98 ;
    END
  END DATA_OUT[0]
  PIN CLOCK
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 34.98 34.98 35.64 35.64 ;
      LAYER Metal6 ;
	RECT 34.98 34.98 35.64 35.64 ;
      LAYER Metal3 ;
	RECT 34.98 34.98 35.64 35.64 ;
      LAYER Metal4 ;
	RECT 34.98 34.98 35.64 35.64 ;
    END
  END CLOCK
  PIN WR_ENABLE
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 42.64 42.64 43.3 43.3 ;
      LAYER Metal6 ;
	RECT 42.64 42.64 43.3 43.3 ;
      LAYER Metal3 ;
	RECT 42.64 42.64 43.3 43.3 ;
      LAYER Metal4 ;
	RECT 42.64 42.64 43.3 43.3 ;
    END
  END WR_ENABLE
  PIN ENABLE
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 50.3 50.3 50.96 50.96 ;
      LAYER Metal6 ;
	RECT 50.3 50.3 50.96 50.96 ;
      LAYER Metal3 ;
	RECT 50.3 50.3 50.96 50.96 ;
      LAYER Metal4 ;
	RECT 50.3 50.3 50.96 50.96 ;
    END
  END ENABLE
    
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 0 70.96 70.96 75.96 ;
        RECT 0 0 70.96 5 ;
      LAYER Metal2 ;
        RECT 65.96 75.96 70.96 5 ;
        RECT 0 0 5 75.96 ;
    END
  END VDD    
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 5.6 62.96 62.96 67.96 ;
        RECT 5.6 5.6 62.96 5 ;
      LAYER Metal2 ;
        RECT 57.96 67.96 62.96 5 ;
        RECT 5.6 5.6 5 67.96 ;
    END
  END VSS    
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 0 78.62 78.62 83.62 ;
        RECT 0 0 78.62 5 ;
      LAYER Metal2 ;
        RECT 73.62 83.62 78.62 5 ;
        RECT 0 0 5 83.62 ;
    END
  END VDD    
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 5.6 70.62 70.62 75.62 ;
        RECT 5.6 5.6 70.62 5 ;
      LAYER Metal2 ;
        RECT 65.62 75.62 70.62 5 ;
        RECT 5.6 5.6 5 75.62 ;
    END
  END VSS