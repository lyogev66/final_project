##
##  Automaticly created by Ofir Even-chen and Yogev Laks Script
####
##  Automaticly created by Ofir Even-chen and Yogev Laks Script
##

VERSION 5.6 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MACRO CDK_R256X16
  CLASS BLOCK ;
  SIZE X_VALUE_SWITCH_LATER BY Y_VALUE_SWITCH_LATER ;
  FOREIGN CDK_R256X16 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN ADDRESS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 12.0 12.0 12.66 12.66 ;
      LAYER Metal6 ;
	RECT 12.0 12.0 12.66 12.66 ;
      LAYER Metal3 ;
	RECT 12.0 12.0 12.66 12.66 ;
      LAYER Metal4 ;
	RECT 12.0 12.0 12.66 12.66 ;
    END
  END ADDRESS[0]
  PIN ADDRESS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 12.0 19.66 12.66 20.32 ;
      LAYER Metal6 ;
	RECT 12.0 19.66 12.66 20.32 ;
      LAYER Metal3 ;
	RECT 12.0 19.66 12.66 20.32 ;
      LAYER Metal4 ;
	RECT 12.0 19.66 12.66 20.32 ;
    END
  END ADDRESS[1]
  PIN ADDRESS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 12.0 27.32 12.66 27.98 ;
      LAYER Metal6 ;
	RECT 12.0 27.32 12.66 27.98 ;
      LAYER Metal3 ;
	RECT 12.0 27.32 12.66 27.98 ;
      LAYER Metal4 ;
	RECT 12.0 27.32 12.66 27.98 ;
    END
  END ADDRESS[2]
  PIN ADDRESS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 12.0 34.98 12.66 35.64 ;
      LAYER Metal6 ;
	RECT 12.0 34.98 12.66 35.64 ;
      LAYER Metal3 ;
	RECT 12.0 34.98 12.66 35.64 ;
      LAYER Metal4 ;
	RECT 12.0 34.98 12.66 35.64 ;
    END
  END ADDRESS[3]
  PIN ADDRESS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 12.0 42.64 12.66 43.3 ;
      LAYER Metal6 ;
	RECT 12.0 42.64 12.66 43.3 ;
      LAYER Metal3 ;
	RECT 12.0 42.64 12.66 43.3 ;
      LAYER Metal4 ;
	RECT 12.0 42.64 12.66 43.3 ;
    END
  END ADDRESS[4]
  PIN ADDRESS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 12.0 50.3 12.66 50.96 ;
      LAYER Metal6 ;
	RECT 12.0 50.3 12.66 50.96 ;
      LAYER Metal3 ;
	RECT 12.0 50.3 12.66 50.96 ;
      LAYER Metal4 ;
	RECT 12.0 50.3 12.66 50.96 ;
    END
  END ADDRESS[5]
  PIN ADDRESS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 12.0 57.96 12.66 58.62 ;
      LAYER Metal6 ;
	RECT 12.0 57.96 12.66 58.62 ;
      LAYER Metal3 ;
	RECT 12.0 57.96 12.66 58.62 ;
      LAYER Metal4 ;
	RECT 12.0 57.96 12.66 58.62 ;
    END
  END ADDRESS[6]
  PIN ADDRESS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 12.0 65.62 12.66 66.28 ;
      LAYER Metal6 ;
	RECT 12.0 65.62 12.66 66.28 ;
      LAYER Metal3 ;
	RECT 12.0 65.62 12.66 66.28 ;
      LAYER Metal4 ;
	RECT 12.0 65.62 12.66 66.28 ;
    END
  END ADDRESS[7]
  PIN DATA_IN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 19.66 12.0 20.32 12.66 ;
      LAYER Metal6 ;
	RECT 19.66 12.0 20.32 12.66 ;
      LAYER Metal3 ;
	RECT 19.66 12.0 20.32 12.66 ;
      LAYER Metal4 ;
	RECT 19.66 12.0 20.32 12.66 ;
    END
  END DATA_IN[0]
  PIN DATA_IN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 27.32 12.0 27.98 12.66 ;
      LAYER Metal6 ;
	RECT 27.32 12.0 27.98 12.66 ;
      LAYER Metal3 ;
	RECT 27.32 12.0 27.98 12.66 ;
      LAYER Metal4 ;
	RECT 27.32 12.0 27.98 12.66 ;
    END
  END DATA_IN[1]
  PIN DATA_IN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 34.98 12.0 35.64 12.66 ;
      LAYER Metal6 ;
	RECT 34.98 12.0 35.64 12.66 ;
      LAYER Metal3 ;
	RECT 34.98 12.0 35.64 12.66 ;
      LAYER Metal4 ;
	RECT 34.98 12.0 35.64 12.66 ;
    END
  END DATA_IN[2]
  PIN DATA_IN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 42.64 12.0 43.3 12.66 ;
      LAYER Metal6 ;
	RECT 42.64 12.0 43.3 12.66 ;
      LAYER Metal3 ;
	RECT 42.64 12.0 43.3 12.66 ;
      LAYER Metal4 ;
	RECT 42.64 12.0 43.3 12.66 ;
    END
  END DATA_IN[3]
  PIN DATA_IN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 50.3 12.0 50.96 12.66 ;
      LAYER Metal6 ;
	RECT 50.3 12.0 50.96 12.66 ;
      LAYER Metal3 ;
	RECT 50.3 12.0 50.96 12.66 ;
      LAYER Metal4 ;
	RECT 50.3 12.0 50.96 12.66 ;
    END
  END DATA_IN[4]
  PIN DATA_IN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 57.96 12.0 58.62 12.66 ;
      LAYER Metal6 ;
	RECT 57.96 12.0 58.62 12.66 ;
      LAYER Metal3 ;
	RECT 57.96 12.0 58.62 12.66 ;
      LAYER Metal4 ;
	RECT 57.96 12.0 58.62 12.66 ;
    END
  END DATA_IN[5]
  PIN DATA_IN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 65.62 12.0 66.28 12.66 ;
      LAYER Metal6 ;
	RECT 65.62 12.0 66.28 12.66 ;
      LAYER Metal3 ;
	RECT 65.62 12.0 66.28 12.66 ;
      LAYER Metal4 ;
	RECT 65.62 12.0 66.28 12.66 ;
    END
  END DATA_IN[6]
  PIN DATA_IN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 73.28 12.0 73.94 12.66 ;
      LAYER Metal6 ;
	RECT 73.28 12.0 73.94 12.66 ;
      LAYER Metal3 ;
	RECT 73.28 12.0 73.94 12.66 ;
      LAYER Metal4 ;
	RECT 73.28 12.0 73.94 12.66 ;
    END
  END DATA_IN[7]
  PIN DATA_IN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 80.94 12.0 81.6 12.66 ;
      LAYER Metal6 ;
	RECT 80.94 12.0 81.6 12.66 ;
      LAYER Metal3 ;
	RECT 80.94 12.0 81.6 12.66 ;
      LAYER Metal4 ;
	RECT 80.94 12.0 81.6 12.66 ;
    END
  END DATA_IN[8]
  PIN DATA_IN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 88.6 12.0 89.26 12.66 ;
      LAYER Metal6 ;
	RECT 88.6 12.0 89.26 12.66 ;
      LAYER Metal3 ;
	RECT 88.6 12.0 89.26 12.66 ;
      LAYER Metal4 ;
	RECT 88.6 12.0 89.26 12.66 ;
    END
  END DATA_IN[9]
  PIN DATA_IN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 96.26 12.0 96.92 12.66 ;
      LAYER Metal6 ;
	RECT 96.26 12.0 96.92 12.66 ;
      LAYER Metal3 ;
	RECT 96.26 12.0 96.92 12.66 ;
      LAYER Metal4 ;
	RECT 96.26 12.0 96.92 12.66 ;
    END
  END DATA_IN[10]
  PIN DATA_IN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 103.92 12.0 104.58 12.66 ;
      LAYER Metal6 ;
	RECT 103.92 12.0 104.58 12.66 ;
      LAYER Metal3 ;
	RECT 103.92 12.0 104.58 12.66 ;
      LAYER Metal4 ;
	RECT 103.92 12.0 104.58 12.66 ;
    END
  END DATA_IN[11]
  PIN DATA_IN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 111.58 12.0 112.24 12.66 ;
      LAYER Metal6 ;
	RECT 111.58 12.0 112.24 12.66 ;
      LAYER Metal3 ;
	RECT 111.58 12.0 112.24 12.66 ;
      LAYER Metal4 ;
	RECT 111.58 12.0 112.24 12.66 ;
    END
  END DATA_IN[12]
  PIN DATA_IN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 119.24 12.0 119.9 12.66 ;
      LAYER Metal6 ;
	RECT 119.24 12.0 119.9 12.66 ;
      LAYER Metal3 ;
	RECT 119.24 12.0 119.9 12.66 ;
      LAYER Metal4 ;
	RECT 119.24 12.0 119.9 12.66 ;
    END
  END DATA_IN[13]
  PIN DATA_IN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 126.9 12.0 127.56 12.66 ;
      LAYER Metal6 ;
	RECT 126.9 12.0 127.56 12.66 ;
      LAYER Metal3 ;
	RECT 126.9 12.0 127.56 12.66 ;
      LAYER Metal4 ;
	RECT 126.9 12.0 127.56 12.66 ;
    END
  END DATA_IN[14]
  PIN DATA_IN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 134.56 12.0 135.22 12.66 ;
      LAYER Metal6 ;
	RECT 134.56 12.0 135.22 12.66 ;
      LAYER Metal3 ;
	RECT 134.56 12.0 135.22 12.66 ;
      LAYER Metal4 ;
	RECT 134.56 12.0 135.22 12.66 ;
    END
  END DATA_IN[15]
  PIN DATA_OUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 142.22 12.0 142.88 12.66 ;
      LAYER Metal6 ;
	RECT 142.22 12.0 142.88 12.66 ;
      LAYER Metal3 ;
	RECT 142.22 12.0 142.88 12.66 ;
      LAYER Metal4 ;
	RECT 142.22 12.0 142.88 12.66 ;
    END
  END DATA_OUT[0]
  PIN DATA_OUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 149.88 12.0 150.54 12.66 ;
      LAYER Metal6 ;
	RECT 149.88 12.0 150.54 12.66 ;
      LAYER Metal3 ;
	RECT 149.88 12.0 150.54 12.66 ;
      LAYER Metal4 ;
	RECT 149.88 12.0 150.54 12.66 ;
    END
  END DATA_OUT[1]
  PIN DATA_OUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 157.54 12.0 158.2 12.66 ;
      LAYER Metal6 ;
	RECT 157.54 12.0 158.2 12.66 ;
      LAYER Metal3 ;
	RECT 157.54 12.0 158.2 12.66 ;
      LAYER Metal4 ;
	RECT 157.54 12.0 158.2 12.66 ;
    END
  END DATA_OUT[2]
  PIN DATA_OUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 165.2 12.0 165.86 12.66 ;
      LAYER Metal6 ;
	RECT 165.2 12.0 165.86 12.66 ;
      LAYER Metal3 ;
	RECT 165.2 12.0 165.86 12.66 ;
      LAYER Metal4 ;
	RECT 165.2 12.0 165.86 12.66 ;
    END
  END DATA_OUT[3]
  PIN DATA_OUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 172.86 12.0 173.52 12.66 ;
      LAYER Metal6 ;
	RECT 172.86 12.0 173.52 12.66 ;
      LAYER Metal3 ;
	RECT 172.86 12.0 173.52 12.66 ;
      LAYER Metal4 ;
	RECT 172.86 12.0 173.52 12.66 ;
    END
  END DATA_OUT[4]
  PIN DATA_OUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 180.52 12.0 181.18 12.66 ;
      LAYER Metal6 ;
	RECT 180.52 12.0 181.18 12.66 ;
      LAYER Metal3 ;
	RECT 180.52 12.0 181.18 12.66 ;
      LAYER Metal4 ;
	RECT 180.52 12.0 181.18 12.66 ;
    END
  END DATA_OUT[5]
  PIN DATA_OUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 188.18 12.0 188.84 12.66 ;
      LAYER Metal6 ;
	RECT 188.18 12.0 188.84 12.66 ;
      LAYER Metal3 ;
	RECT 188.18 12.0 188.84 12.66 ;
      LAYER Metal4 ;
	RECT 188.18 12.0 188.84 12.66 ;
    END
  END DATA_OUT[6]
  PIN DATA_OUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 195.84 12.0 196.5 12.66 ;
      LAYER Metal6 ;
	RECT 195.84 12.0 196.5 12.66 ;
      LAYER Metal3 ;
	RECT 195.84 12.0 196.5 12.66 ;
      LAYER Metal4 ;
	RECT 195.84 12.0 196.5 12.66 ;
    END
  END DATA_OUT[7]
  PIN DATA_OUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 203.5 12.0 204.16 12.66 ;
      LAYER Metal6 ;
	RECT 203.5 12.0 204.16 12.66 ;
      LAYER Metal3 ;
	RECT 203.5 12.0 204.16 12.66 ;
      LAYER Metal4 ;
	RECT 203.5 12.0 204.16 12.66 ;
    END
  END DATA_OUT[8]
  PIN DATA_OUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 211.16 12.0 211.82 12.66 ;
      LAYER Metal6 ;
	RECT 211.16 12.0 211.82 12.66 ;
      LAYER Metal3 ;
	RECT 211.16 12.0 211.82 12.66 ;
      LAYER Metal4 ;
	RECT 211.16 12.0 211.82 12.66 ;
    END
  END DATA_OUT[9]
  PIN DATA_OUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 218.82 12.0 219.48 12.66 ;
      LAYER Metal6 ;
	RECT 218.82 12.0 219.48 12.66 ;
      LAYER Metal3 ;
	RECT 218.82 12.0 219.48 12.66 ;
      LAYER Metal4 ;
	RECT 218.82 12.0 219.48 12.66 ;
    END
  END DATA_OUT[10]
  PIN DATA_OUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 226.48 12.0 227.14 12.66 ;
      LAYER Metal6 ;
	RECT 226.48 12.0 227.14 12.66 ;
      LAYER Metal3 ;
	RECT 226.48 12.0 227.14 12.66 ;
      LAYER Metal4 ;
	RECT 226.48 12.0 227.14 12.66 ;
    END
  END DATA_OUT[11]
  PIN DATA_OUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 234.14 12.0 234.8 12.66 ;
      LAYER Metal6 ;
	RECT 234.14 12.0 234.8 12.66 ;
      LAYER Metal3 ;
	RECT 234.14 12.0 234.8 12.66 ;
      LAYER Metal4 ;
	RECT 234.14 12.0 234.8 12.66 ;
    END
  END DATA_OUT[12]
  PIN DATA_OUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 241.8 12.0 242.46 12.66 ;
      LAYER Metal6 ;
	RECT 241.8 12.0 242.46 12.66 ;
      LAYER Metal3 ;
	RECT 241.8 12.0 242.46 12.66 ;
      LAYER Metal4 ;
	RECT 241.8 12.0 242.46 12.66 ;
    END
  END DATA_OUT[13]
  PIN DATA_OUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 249.46 12.0 250.12 12.66 ;
      LAYER Metal6 ;
	RECT 249.46 12.0 250.12 12.66 ;
      LAYER Metal3 ;
	RECT 249.46 12.0 250.12 12.66 ;
      LAYER Metal4 ;
	RECT 249.46 12.0 250.12 12.66 ;
    END
  END DATA_OUT[14]
  PIN DATA_OUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 257.12 12.0 257.78 12.66 ;
      LAYER Metal6 ;
	RECT 257.12 12.0 257.78 12.66 ;
      LAYER Metal3 ;
	RECT 257.12 12.0 257.78 12.66 ;
      LAYER Metal4 ;
	RECT 257.12 12.0 257.78 12.66 ;
    END
  END DATA_OUT[15]
  PIN CLOCK
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 264.78 12.0 265.44 12.66 ;
      LAYER Metal6 ;
	RECT 264.78 12.0 265.44 12.66 ;
      LAYER Metal3 ;
	RECT 264.78 12.0 265.44 12.66 ;
      LAYER Metal4 ;
	RECT 264.78 12.0 265.44 12.66 ;
    END
  END CLOCK
  PIN WR_ENABLE
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 272.44 12.0 273.1 12.66 ;
      LAYER Metal6 ;
	RECT 272.44 12.0 273.1 12.66 ;
      LAYER Metal3 ;
	RECT 272.44 12.0 273.1 12.66 ;
      LAYER Metal4 ;
	RECT 272.44 12.0 273.1 12.66 ;
    END
  END WR_ENABLE
  PIN ENABLE
    DIRECTION INPUT ;
    USE SIGNAL ;
  PORT
      LAYER Metal5 ;
	RECT 280.1 12.0 280.76 12.66 ;
      LAYER Metal6 ;
	RECT 280.1 12.0 280.76 12.66 ;
      LAYER Metal3 ;
	RECT 280.1 12.0 280.76 12.66 ;
      LAYER Metal4 ;
	RECT 280.1 12.0 280.76 12.66 ;
    END
  END ENABLE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 0 79.28 293.76 84.28 ;
        RECT 0 0 293.76 5 ;
      LAYER Metal2 ;
        RECT 288.76 84.28 293.76 5 ;
        RECT 0 0 5 84.28 ;
    END
  END VDD    
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 5.6 71.28 285.76 76.28 ;
        RECT 5.6 5.6 285.76 5 ;
      LAYER Metal2 ;
        RECT 280.76 76.28 285.76 5 ;
        RECT 5.6 5.6 5 76.28 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 12.0 12.0 280.76 66.28 ;
    LAYER Metal2 ;
      RECT 12.0 12.0 280.76 66.28 ;
    LAYER Metal3 ;
      RECT 12.0 12.0 280.76 66.28 ;
    LAYER Metal4 ;
      RECT 12.0 12.0 280.76 66.28 ;
    LAYER Metal5 ;
      RECT 12.0 12.0 280.76 66.28 ;
    LAYER Metal6 ;
      RECT 12.0 12.0 280.76 66.28 ;
  END
END CDK_R512x16

END LIBRARY
    